;HorizontalDatum:  UTMNAD83
;HorizontalZone:   10
;HorizontalUnits:  Meters
;VerticalDatum:    NAVD88
;VerticalUnits:    USSurveyFeet
;Filetype:          landmark
;NumElements:      432
586698.56,4214178.0,329
594099.1,4214269.0,328
587744.0,4223991.5,327
611430.2,4235208.0,326
609135.1,4235300.5,325
607129.5,4235391.5,324
615267.7,4233075.5,323
614731.2,4233715.5,322
614325.75,4235208.0,321
627840.56,4231551.5,289
611582.6,4238622.5,320
628919.56,4231855.5,288
626240.3,4222376.5,287
627569.25,4223108.5,286
628788.44,4225515.5,285
628928.6,4226857.5,284
629145.06,4228746.5,283
630391.6,4229417.5,282
630928.06,4230301.5,281
630760.5,4231733.5,280
614182.56,4243133.5,319
616746.0,4238622.5,318
616483.75,4243895.5,317
616017.5,4232160.0,316
616992.75,4236793.5,315
618262.25,4244148.5,314
619714.7,4248802.5,313
621997.7,4254776.0,312
623488.06,4259165.0,311
634533.8,4222407.5,279
623344.94,4266572.0,310
637508.6,4223229.5,278
634454.56,4225637.5,277
635564.06,4229569.5,275
605245.75,4236976.5,273
624347.5,4219023.5,272
624816.94,4221157.5,271
626871.2,4219755.5,270
628051.06,4269071.0,309
618934.3,4236519.5,308
618431.5,4238744.0,307
620622.94,4228137.5,306
622308.5,4232221.5,305
622421.25,4234873.5,304
623268.6,4237342.5,303
621945.7,4238439.5,302
629266.9,4220334.5,269
622720.0,4241243.5,301
631699.1,4219724.5,268
623753.2,4243560.5,300
631296.8,4221157.5,267
631016.5,4222285.5,266
631104.9,4223473.5,265
632046.7,4225150.5,264
632269.2,4226948.5,263
633180.56,4228411.5,262
631891.4,4230301.5,261
631909.6,4232099.5,260
632592.3,4233623.5,259
633326.94,4235391.5,258
636551.75,4235269.0,257
631385.4,4233014.5,256
631537.75,4233715.5,255
631351.9,4235086.5,254
631549.94,4236214.5,253
627462.5,4216463.5,252
629827.75,4216585.5,251
632122.8,4217042.5,250
632217.4,4218505.5,249
634110.1,4216189.5,248
635176.94,4214482.5,247
638861.94,4216493.5,246
631345.6,4214756.5,245
633384.7,4211434.5,244
635158.56,4212775.5,243
638636.4,4211799.5,242
641879.4,4208477.5,241
615395.7,4219328.5,240
620171.75,4219633.5,239
588070.25,4215427.5,238
612320.2,4208387.0,237
615517.44,4208173.0,236
622424.2,4211709.0,235
621299.5,4210977.5,234
624155.4,4211709.0,232
622326.56,4198755.0,199
623853.7,4213080.5,231
622521.7,4197535.5,198
621174.5,4212775.5,230
624021.25,4197870.5,197
625121.6,4197658.0,196
627492.94,4197139.5,195
628977.3,4197170.0,194
623765.3,4188117.5,193
627304.0,4191378.5,192
628837.1,4192292.8,191
629663.1,4192749.5,190
590536.06,4213750.5,227
618586.75,4212805.5,226
620177.9,4212197.0,225
622524.9,4213415.5,224
615450.44,4208326.0,223
618958.56,4208112.0,222
630522.6,4193207.8,189
616431.9,4210001.5,221
631924.75,4193999.5,188
618211.9,4211860.5,220
627691.0,4190677.5,187
628358.44,4190951.5,186
628321.94,4190159.8,185
628940.75,4190098.8,184
628748.75,4189549.8,183
628343.3,4188513.8,182
624569.94,4184215.8,181
625085.0,4185831.5,180
621284.2,4210215.5,219
620385.06,4207625.0,218
621445.8,4207899.0,217
622280.9,4208630.5,216
620884.9,4206314.0,215
620970.3,4204516.0,214
627489.9,4200095.5,213
624923.44,4191286.5,212
625460.0,4186288.8,179
624463.25,4189945.8,211
628824.94,4186745.8,178
623868.8,4189153.5,210
630894.5,4186775.8,177
632150.2,4186806.5,176
633326.8,4186836.8,175
634356.94,4186836.8,174
635673.75,4186867.5,173
636444.94,4186897.8,172
638227.94,4186958.8,171
640318.9,4186989.8,170
622945.3,4188757.8,209
627032.75,4207899.0,208
628669.4,4207350.0,207
619367.0,4203997.5,206
620970.3,4204210.5,205
622558.3,4204089.0,204
623472.6,4203570.5,203
622686.3,4202686.5,202
639538.6,4185160.8,169
622305.3,4201558.5,201
641525.9,4185404.2,168
622134.56,4199912.5,200
643501.0,4184703.5,167
645314.6,4183209.2,166
643501.0,4185038.5,165
645354.25,4183819.2,164
646829.44,4182142.2,163
648865.5,4180466.5,162
639547.75,4183057.5,160
640008.0,4182417.8,159
641373.5,4181838.8,157
641931.3,4182264.8,156
642208.56,4181533.5,155
642979.8,4181259.2,154
639285.6,4183666.5,149
634488.06,4202808.5,148
635920.56,4201833.5,147
637810.4,4199729.5,146
629794.06,4203631.5,145
631110.9,4203661.5,144
632397.06,4203661.5,143
633945.44,4203692.5,142
634030.8,4205002.5,141
635487.7,4205825.5,140
642345.75,4202381.5,139
643007.1,4200888.5,138
631156.56,4206130.5,137
630562.2,4205460.5,136
630394.56,4204516.0,135
629163.2,4211556.5,134
630138.56,4209178.5,133
630187.25,4207929.5,132
630870.06,4207868.5,131
630653.7,4207076.0,130
629855.06,4206984.5,129
629111.4,4206191.5,128
628727.3,4205307.5,127
628706.0,4204363.0,126
628718.25,4203387.5,125
629080.94,4202168.5,124
629608.25,4201041.0,123
628733.44,4200980.0,122
628876.75,4200065.5,121
629373.5,4199303.5,120
629303.44,4198267.0,119
630132.5,4197932.0,118
630464.75,4197352.5,117
631101.75,4196529.5,116
631973.44,4196224.5,115
632256.9,4195523.5,114
632851.25,4194517.5,113
634689.2,4193847.8,112
636652.06,4194243.8,111
637859.06,4195005.5,110
639291.6,4194578.5,109
641038.1,4194395.5,108
642178.2,4193329.2,107
642818.25,4191530.5,106
642574.44,4190159.5,105
641995.3,4188025.5,104
624402.3,4213537.5,103
624560.8,4210245.5,102
624976.56,4211592.5,101
626657.75,4208691.5,100
624676.5,4207441.5,99
625645.8,4206831.5,98
624716.25,4206435.5,97
625130.8,4206040.0,96
624646.1,4205490.5,95
624579.0,4204759.5,94
625051.56,4203754.0,93
625392.8,4202747.5,92
626075.6,4202230.0,91
625176.5,4201742.0,90
630662.94,4235818.5,455
631470.6,4236915.5,454
630699.56,4238988.5,453
630166.2,4240999.0,452
631199.5,4242462.0,451
630888.6,4243072.0,450
626222.0,4201619.5,89
625780.0,4200553.0,88
626718.7,4200796.5,87
626468.8,4200095.5,86
626822.3,4199120.5,85
626999.1,4198083.5,84
626081.75,4197413.5,83
634442.44,4236854.0,449
626292.06,4197078.5,82
636405.44,4238134.0,448
625487.3,4196041.5,81
637249.6,4235208.0,447
625999.44,4195005.5,80
637130.8,4235482.0,446
581364.56,4223535.0,445
579221.8,4219360.0,444
579925.9,4223017.0,443
578840.8,4220274.0,442
579782.7,4218933.0,440
625237.44,4194273.5,79
625103.3,4193024.5,78
625490.44,4191835.8,77
625907.94,4191256.8,76
626429.2,4190707.8,75
626758.3,4189671.8,74
627044.8,4188787.8,73
627386.25,4187812.8,72
579791.8,4220152.0,438
627474.7,4187355.5,71
626929.0,4186410.8,70
588570.0,4218018.0,436
591517.56,4216920.5,434
593818.75,4216585.5,433
586671.06,4226521.5,399
585040.5,4227527.5,398
585046.6,4228929.5,397
578139.8,4231064.0,396
586180.4,4231276.5,395
582788.06,4228563.5,394
581358.56,4228807.5,393
583095.9,4231460.0,392
578414.06,4224907.0,391
580322.2,4226583.0,390
628261.0,4185709.8,69
629120.5,4185129.5,68
629855.1,4184398.8,67
631400.44,4183453.8,66
632348.44,4182600.8,65
633409.1,4182691.8,64
634158.94,4183453.8,63
634820.3,4184459.8,62
583086.7,4223383.0,428
635719.5,4184947.8,61
637060.6,4184916.5,60
588518.2,4226675.0,425
591301.06,4225333.5,422
593355.44,4224845.5,421
578938.4,4226827.0,389
595611.0,4221949.5,420
581285.4,4226157.0,388
581431.6,4227344.5,387
579730.8,4223901.0,386
578725.0,4215824.0,385
578981.0,4218598.0,384
579237.06,4221463.0,383
578688.4,4223718.0,382
577819.7,4224694.0,381
577771.0,4227802.0,380
637813.4,4184428.5,59
639087.44,4184672.8,58
639050.94,4185160.8,57
639191.1,4186013.8,56
641656.94,4185861.5,54
642598.8,4186989.5,53
643019.44,4187233.2,52
597747.7,4216432.5,418
644314.8,4186928.2,51
597976.3,4214847.5,417
645366.4,4187263.5,50
597918.44,4215579.5,415
591672.94,4226704.5,413
595696.44,4225425.0,412
576527.4,4229448.0,379
595559.2,4226461.0,410
581096.3,4219695.0,378
580389.2,4221249.0,377
582553.4,4223718.0,376
582056.5,4225242.0,375
583318.4,4226034.5,374
584205.3,4227527.5,373
584357.75,4229752.5,372
584851.56,4230606.5,371
575783.7,4230210.0,370
646070.5,4187294.2,49
541536.6,4184108.0,806
646515.5,4186410.2,48
546104.3,4185736.5,805
602627.5,4209666.5,47
550155.7,4193402.0,804
606937.44,4208508.5,46
548924.4,4200750.0,803
611594.7,4209940.5,45
549718.75,4203967.0,802
615700.44,4213323.5,44
558536.4,4211593.5,801
615621.1,4215914.5,43
564719.56,4212888.0,800
594775.94,4228503.5,409
618888.56,4216432.5,42
596418.7,4231093.5,408
621476.25,4218078.5,41
624917.4,4217133.5,40
594720.94,4226126.0,406
587356.94,4231276.5,405
588545.7,4231154.5,404
593855.4,4230087.5,403
584589.44,4226217.5,402
586393.8,4226247.5,401
575244.2,4230363.0,369
584702.1,4218841.0,368
579898.5,4214940.0,367
584113.94,4215092.0,366
582632.5,4218872.0,365
582745.3,4220457.0,364
585650.06,4216982.0,363
588499.94,4212562.0,362
575853.8,4209728.0,361
577182.7,4210734.0,360
625127.8,4216097.5,39
625621.5,4215030.5,38
627054.06,4213202.5,37
628660.3,4214299.5,36
628608.5,4212958.5,35
630028.8,4212744.5,34
631497.4,4211860.5,33
632622.7,4210977.5,32
632400.2,4210154.5,31
634128.4,4209879.5,30
581023.2,4212380.0,359
585644.0,4213142.0,358
592300.9,4212714.5,357
597549.5,4211556.5,356
601076.1,4214055.5,355
605187.8,4212988.5,354
610418.25,4216250.5,353
613332.1,4218718.5,352
614844.0,4222528.5,351
616736.7,4226277.5,350
635371.94,4208416.5,29
635079.4,4207380.5,28
636764.9,4207959.5,27
636630.7,4206618.5,26
637517.7,4206191.5,25
639508.06,4206252.0,24
640471.2,4205764.5,23
641995.2,4204667.5,22
643214.44,4203326.5,21
644137.9,4202473.5,20
619586.6,4225698.5,349
622043.25,4224875.5,348
648365.6,4187690.2,9
624067.06,4227314.0,347
647228.7,4185800.5,8
626270.9,4229112.0,346
648490.56,4184093.2,7
626273.9,4231002.5,345
649615.3,4182600.2,6
626301.3,4233288.5,344
649395.75,4179704.5,5
629763.9,4233440.5,343
649947.44,4176687.2,4
630306.4,4234233.5,342
651800.7,4176016.5,3
627682.1,4237250.5,341
652401.25,4174797.5,2
624743.8,4240573.5,340
651986.6,4172328.2,1
645098.0,4202046.5,19
646201.4,4201650.5,18
645793.0,4201131.5,17
645320.7,4200644.0,16
646280.7,4200187.5,15
646932.9,4199181.5,14
647716.3,4198266.5,13
646942.1,4195279.5,12
647509.06,4192048.2,11
647472.4,4190098.5,10
624527.5,4243072.5,339
628264.2,4245937.0,338
629187.8,4249229.0,337
628383.1,4253892.0,336
630623.5,4255721.0,335
628532.56,4259409.0,334
625633.9,4262152.0,333
628624.0,4264591.0,332
628910.56,4269163.0,331
624725.5,4246059.0,299
629904.3,4272881.0,330
626420.2,4247888.0,298
627633.4,4250326.0,297
628739.7,4252643.0,296
623158.75,4221797.5,295
623780.56,4223016.0,294
624082.4,4224936.5,293
624969.4,4226887.5,292
626852.94,4228228.5,291
628172.75,4230209.5,290
